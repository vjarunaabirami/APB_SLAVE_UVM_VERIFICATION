
`include "uvm_macros.svh"
package apb_slave_package;
import uvm_pkg::*;
//`include "uvm_macros.svh"
`include "defines.sv"
`include "apb_slave_sequence_item.sv"
`include "apb_slave_sequence.sv"
`include "apb_slave_sequencer.sv"
`include "apb_slave_driver.sv"
`include "apb_slave_active_monitor.sv"
`include "apb_slave_passive_monitor.sv"
`include "apb_slave_active_agent.sv"
`include "apb_slave_passive_agent.sv"
`include "apb_slave_scoreboard.sv"
`include "apb_slave_subscriber.sv"
`include "apb_slave_environment.sv"
`include "apb_slave_test.sv"

endpackage

