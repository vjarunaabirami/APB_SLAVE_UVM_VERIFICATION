 `define ADDR_WIDTH 8
`define DATA_WIDTH 256
`define MEM_DEPTH  256
